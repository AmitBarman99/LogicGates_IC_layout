*** SPICE deck for cell NOR{lay} from library NORgate
*** Created on Thu Jul 07, 2022 23:29:46
*** Last revised on Fri Jul 08, 2022 01:31:30
*** Written on Fri Jul 08, 2022 01:33:15 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NOR{lay}
Mnmos@0 gnd net@15 AnorB gnd NMOS L=0.36U W=1.8U AS=1.944P AD=5.184P PS=4.56U PD=13.32U
Mnmos@1 AnorB A gnd gnd NMOS L=0.36U W=1.8U AS=5.184P AD=1.944P PS=13.32U PD=4.56U
Mpmos@0 vdd net@15 net@11 vdd PMOS L=0.36U W=1.8U AS=0.972P AD=9.007P PS=2.88U PD=20.52U
Mpmos@1 net@11 A AnorB vdd PMOS L=0.36U W=1.8U AS=1.944P AD=0.972P PS=4.56U PD=2.88U

* Spice Code nodes in cell cell 'NOR{lay}'
vdd vdd 0 DC 5
va A 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb B 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.measure tran tf trig v(AnorB) val=4.5 fall=1 td=4ns trag v(AnorB) val=0.5 fall=1
.measure tran tr trig v(AnorB) val=0.5 rise=1 td=4ns trag v(AnorB) val=4.5 rise=1
.tran 200n
.include D:\Electric\projects\C5_models.txt
.END
